library verilog;
use verilog.vl_types.all;
entity tristate_driver_tb is
end tristate_driver_tb;
