library verilog;
use verilog.vl_types.all;
entity bitwise_comparator_tb is
end bitwise_comparator_tb;
