library verilog;
use verilog.vl_types.all;
entity bitwise_and_tb is
end bitwise_and_tb;
