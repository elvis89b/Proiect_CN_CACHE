library verilog;
use verilog.vl_types.all;
entity bit_comparator_tb is
end bit_comparator_tb;
