module cache_controller #(parameter ADDRESS_WORD_SIZE = 32, parameter TAG_SIZE = 19, parameter BLOCK_SIZE = 8, parameter WORD_SIZE = 8, parameter NUMBER_OF_SETS = 128) (
  input clk,
  input rst_b,
  input opcode, // 1 - write, 0 - read
  output [7:0]data,
  output hit_miss
);

  // internal wires
  wire hit_miss_w;
  wire [3:0]hit_miss_set;
  wire [7:0]ages;
  wire [ADDRESS_WORD_SIZE-1:0]address_word;
  wire try_read;
  wire try_write;
  wire [7:0]write_data;
  wire [3:0]reset_age;
  wire [3:0]increment_age;
  
  
  // instantiate the control unit
  control_unit #(.ADDRESS_WORD_SIZE(ADDRESS_WORD_SIZE)) uut_control (
    .clk(clk),
    .rst_b(rst_b),
    .opcode(opcode),
    .hit_miss(hit_miss_w),
    .hit_miss_set(hit_miss_set),
    .ages(ages),
    .address_word(address_word),
    .try_read(try_read),
    .try_write(try_write),
    .write_data(write_data),
    .reset_age(reset_age),
    .increment_age(increment_age)
  );
  
  // instantiate the cache memory
  cache_memory #(
    .ADDRESS_WORD_SIZE(ADDRESS_WORD_SIZE),
    .TAG_SIZE(TAG_SIZE),
    .BLOCK_SIZE(BLOCK_SIZE),
    .WORD_SIZE(WORD_SIZE),
    .NUMBER_OF_SETS(NUMBER_OF_SETS)
  ) uut_cache (
    .clk(clk),
    .rst_b(rst_b),
    .address_word(address_word),
    .try_read(try_read),
    .try_write(try_write),
    .write_data(write_data),
    .reset_age(reset_age),
    .increment_age(increment_age),
    .data(data),
    .ages(ages),
    .hit_miss(hit_miss_w),
    .hit_miss_set(hit_miss_set)
  );
  
  // send hit_miss signal to output
  assign hit_miss = hit_miss_w;
  
endmodule