library verilog;
use verilog.vl_types.all;
entity mux128to1_tb is
end mux128to1_tb;
