library verilog;
use verilog.vl_types.all;
entity four_way_set_tb is
end four_way_set_tb;
