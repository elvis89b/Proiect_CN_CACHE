library verilog;
use verilog.vl_types.all;
entity cache_line_tb is
end cache_line_tb;
