library verilog;
use verilog.vl_types.all;
entity cache_controller_tb is
end cache_controller_tb;
