library verilog;
use verilog.vl_types.all;
entity cache_memory_tb is
end cache_memory_tb;
