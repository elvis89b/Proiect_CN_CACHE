module bitwise_and (
  input in_0,
  input in_1,
  output and_
);

  assign and_ = in_0 & in_1;
  
endmodule