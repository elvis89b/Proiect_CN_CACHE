library verilog;
use verilog.vl_types.all;
entity dec7to128_tb is
end dec7to128_tb;
