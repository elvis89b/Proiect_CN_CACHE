library verilog;
use verilog.vl_types.all;
entity encoder4to2_tb is
end encoder4to2_tb;
