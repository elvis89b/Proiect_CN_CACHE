library verilog;
use verilog.vl_types.all;
entity and_wordgate_tb is
end and_wordgate_tb;
